`include control.v 
`include ALU.v

module processor();
reg clk;
